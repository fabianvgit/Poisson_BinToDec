library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package data1_types is

type integer_vector is array (natural range <>) of integer;
end data1_types;